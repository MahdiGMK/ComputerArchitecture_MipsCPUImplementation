library verilog;
use verilog.vl_types.all;
entity PipelineCPU_vlg_vec_tst is
end PipelineCPU_vlg_vec_tst;
