library verilog;
use verilog.vl_types.all;
entity Instruction_Memory_vlg_vec_tst is
end Instruction_Memory_vlg_vec_tst;
